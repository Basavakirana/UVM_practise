class rd_agt_config extends uvm_object;

    `uvm_object_utils(rd_agt_config)

    uvm_active_passive_enum is_active = UVM_ACTIVE;

    function new(string name="rd_agt_config");
        super.new(name);
    endfunction
      
endclass

  //  extern function new(string name="rd_agt_config");
