package apb_test_pkg;
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "../uvm_testbench/apb_sequence/apb_seq_item.sv"
`include "../uvm_testbench/apb_sequence/apb_seq_item_slave.sv"
`include "../uvm_testbench/apb_sequence/apb_sequence_slave_rw.sv"
`include "../uvm_testbench/apb_sequence/apb_sequence_write.sv"

`include "../uvm_testbench/apb_agent/apb_sequencer.sv"
`include "../uvm_testbench/apb_agent/apb_driver.sv"
`include "../uvm_testbench/apb_agent/apb_slave_sequencer.sv"
`include "../uvm_testbench/apb_agent/apb_driver_slave.sv"
`include "../uvm_testbench/apb_agent/apb_monitor.sv"
`include "../uvm_testbench/apb_agent/apb_agent_jtag.sv"
`include "../uvm_testbench/apb_agent/apb_agent_slave.sv"

`include "../uvm_testbench/apb_env/apb_scoreboard.sv"
`include "../uvm_testbench/apb_env/apb_env.sv"

`include "../uvm_testbench/apb_test/apb_test.sv"

endpackage

